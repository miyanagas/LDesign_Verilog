module jk_ff (Clk, J, K);
    input Clk, J, K;
    output Q;
    reg Q;

    always @(posedge Clk) begin
        if (J == 1'b1 and K == 1'b1) begin
            Q <= ~Q;
        end
        else if (J | K == 1'b1) begin
            Q <= J;
        end
    end
endmodule